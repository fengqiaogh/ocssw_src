netcdf PACE_OCI.20220321T000000.L1B.rhot-ocean {
dimensions:
	number_of_scans = UNLIMITED ;
//	CCD_pixels = 1272 ;
//	SWIR_pixels = 1272 ;
//	blue_bands = 120 ;
//	red_bands = 120 ;
	SWIR_bands = 9 ;
	vector_elements = 3 ;
	quaternion_elements = 4 ;
	polarization_coefficients = 3 ;
	HAM_sides = 2 ;

// global attributes:
		:title = "PACE OCI Level-1B Data" ;
		:instrument = "OCI" ;
		:date_created = "2022-01-10T10:39:18Z" ;
		:product_name = "PACE_OCI.20190321T062500.L1B.nc" ;
		:processing_version = "V1.0" ;
		:Conventions = "CF-1.8 ACDD-1.3" ;
		:institution = "NASA Goddard Space Flight Center, Ocean Biology Processing Group" ;
		:license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/" ;
		:naming_authority = "gov.nasa.gsfc.oceancolor" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "CF Standard Name Table v79" ;
		:creator_name = "NASA/GSFC/OBPG" ;
		:creator_email = "data@oceancolor.gsfc.nasa.gov" ;
		:creator_url = "https://oceancolor.gsfc.nasa.gov" ;
		:project = "Ocean Biology Processing Group" ;
		:publisher_name = "NASA/GSFC/OB.DAAC" ;
		:publisher_email = "data@oceancolor.gsfc.nasa.gov" ;
		:publisher_url = "https://oceancolor.gsfc.nasa.gov" ;
		:processing_level = "L1B" ;
		:cdm_data_type = "swath" ;
		:normalizedLt = 0 ;
		:sample_offset = 0 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_min = "73.55669f ;" ;
		:geospatial_lat_max = "45.88998f ;" ;
		:geospatial_lon_min = "35.87455f ;" ;
		:geospatial_lon_max = "8.31627f ;" ;
  		:gringpointlongitude = 22.58846f, -5.335992f, -9.173955f, -9.461103f ;
  		:gringpointlatitude = -13.02491f, -17.24885f, 2.346621f, 3.552641f ;
  		:gringpointsequence = 1, 2, 3, 4 ;
		:time_coverage_start = "2019-03-21T06:25:00" ;
		:time_coverage_end = "2019-03-21T06:30:00" ;
		:history = "l1bgeogen_oci" ;
		:earth_sun_distance_correction = 1.00780784057772 ;
		:CDL_version_date = "2024-10-14" ;

group: sensor_band_parameters {
  variables:
//  	float blue_wavelength(blue_bands) ;
//  		blue_wavelength:_FillValue = -32767.f ;
//  		blue_wavelength:long_name = "Band center wavelengths for bands from blue CCD" ;
//  		blue_wavelength:valid_min = 310.f ;
//  		blue_wavelength:valid_max = 610.f ;
//  		blue_wavelength:units = "nm" ;
//  	float red_wavelength(red_bands) ;
//  		red_wavelength:_FillValue = -32767.f ;
//  		red_wavelength:long_name = "Band center wavelengths for bands from red CCD" ;
//  		red_wavelength:valid_min = 595.f ;
//  		red_wavelength:valid_max = 900.f ;
//  		red_wavelength:units = "nm" ;
  	float SWIR_wavelength(SWIR_bands) ;
  		SWIR_wavelength:_FillValue = -32767.f ;
  		SWIR_wavelength:long_name = "Band center wavelengths for SWIR bands" ;
  		SWIR_wavelength:valid_min = 939.f ;
  		SWIR_wavelength:valid_max = 2260.f ;
  		SWIR_wavelength:units = "nm" ;
  	float SWIR_bandpass(SWIR_bands) ;
  		SWIR_bandpass:_FillValue = -32767.f ;
  		SWIR_bandpass:long_name = "Bandpasses for SWIR bands" ;
  		SWIR_bandpass:valid_min = 0.f ;
  		SWIR_bandpass:valid_max = 100.f ;
  		SWIR_bandpass:units = "nm" ;
//  	float blue_solar_irradiance(blue_bands) ;
//  		blue_solar_irradiance:_FillValue = -32767.f ;
//  		blue_solar_irradiance:long_name = "Mean extraterrestrial solar irradiance at 1 astronomical unit for the wavelengths of the blue CCD" ;
//  		blue_solar_irradiance:valid_min = 0.f ;
//  		blue_solar_irradiance:valid_max = 2500.f ;
//  		blue_solar_irradiance:units = "W m^-2 um^-1" ;
//  	float red_solar_irradiance(red_bands) ;
//  		red_solar_irradiance:_FillValue = -32767.f ;
//  		red_solar_irradiance:long_name = "Mean extraterrestrial solar irradiance at 1 astronomical unit for the wavelengths of the red CCD" ;
//  		red_solar_irradiance:valid_min = 0.f ;
//  		red_solar_irradiance:valid_max = 2500.f ;
//  		red_solar_irradiance:units = "W m^-2 um^-1" ;
  	float SWIR_solar_irradiance(SWIR_bands) ;
  		SWIR_solar_irradiance:_FillValue = -32767.f ;
  		SWIR_solar_irradiance:long_name = "Mean extraterrestrial solar irradiance at 1 astronomical unit for the SWIR wavelengths" ;
  		SWIR_solar_irradiance:valid_min = 7.f ;
  		SWIR_solar_irradiance:valid_max = 95.f ;
  		SWIR_solar_irradiance:units = "W m^-2 um^-1" ;
//  	float blue_m12_coef(blue_bands, HAM_sides, polarization_coefficients) ;
//  		blue_m12_coef:long_name = "Blue band M12/M11 polynomial coefficients" ;
//  		blue_m12_coef:units = "dimensionless" ;
//  	float blue_m13_coef(blue_bands, HAM_sides, polarization_coefficients) ;
//  		blue_m13_coef:long_name = "Blue band M13/M11 polynomial coefficients" ;
//  		blue_m13_coef:units = "dimensionless" ;
//  	float red_m12_coef(red_bands, HAM_sides, polarization_coefficients) ;
//  		red_m12_coef:long_name = "Red band m12/M11 polynomial coefficients" ;
//  		red_m12_coef:units = "dimensionless" ;
//  	float red_m13_coef(red_bands, HAM_sides, polarization_coefficients) ;
//  		red_m13_coef:long_name = "Red band M13/M11 polynomial coefficients" ;
//  		red_m13_coef:units = "dimensionless" ;
  	float SWIR_m12_coef(SWIR_bands, HAM_sides, polarization_coefficients) ;
     		SWIR_m12_coef:long_name = "SWIR band M12/M11 polynomial coefficients" ;
  		SWIR_m12_coef:units = "dimensionless" ;
  	float SWIR_m13_coef(SWIR_bands, HAM_sides, polarization_coefficients) ;
  		SWIR_m13_coef:long_name = "SWIR band M13/M11 polynomial coefficients" ;
  		SWIR_m13_coef:units = "dimensionless" ;
  } // group sensor_band_parameters

group: scan_line_attributes {
  variables:
  	double time(number_of_scans) ;
  		time:_FillValue = -32767. ;
  		time:long_name = "time" ;
  		time:units = "seconds since 2022-03-21 00:00:00" ;
  		time:description = "Earth view mid time in seconds of day" ;
  		time:valid_min = 0. ;
  		time:valid_max = 86401. ;
  	ubyte HAM_side(number_of_scans) ;
  		HAM_side:_FillValue = 255UB ;
  		HAM_side:long_name = "Half-angle mirror side" ;
  		HAM_side:valid_min = 0UB ;
  		HAM_side:valid_max = 1UB ;
  	ubyte scan_quality_flags(number_of_scans) ;
  		scan_quality_flags:_FillValue = 255UB ;
  		scan_quality_flags:long_name = "Scan quality flags " ;
  		scan_quality_flags:units = "none" ;
  		scan_quality_flags:flag_masks = 1, 2, 4 ;
  		scan_quality_flags:flag_meanings = "tilt_change missing_time missing_encoder" ;
  } // group scan_line_attributes

//group: geolocation_data {
//  variables:
//  	float latitude(number_of_scans, CCD_pixels) ;
//  		latitude:_FillValue = -32767.f ;
// 		latitude:long_name = "Latitudes of pixel locations" ;
//  		latitude:units = "degrees_north" ;
//		latitude:valid_min = -90.f ;
//		latitude:valid_max = 90.f ;
//	float longitude(number_of_scans, CCD_pixels) ;
//		longitude:_FillValue = -32767.f ;
//		longitude:long_name = "Longitudes of pixel locations" ;
//		longitude:units = "degrees_east" ;
//		longitude:valid_min = -180.f ;
//		longitude:valid_max = 180.f ;
//	short height(number_of_scans, CCD_pixels) ;
//		height:_FillValue = -32767s ;
//		height:long_name = "Terrain height at pixel locations" ;
//		height:units = "meters" ;
//		height:valid_min = -1000s ;
//		height:valid_max = 10000s ;
//		height:scale_factor = 1. ;
//		height:add_offset = 0. ;
//	short sensor_azimuth(number_of_scans, CCD_pixels) ;
//		sensor_azimuth:_FillValue = -32767s ;
//		sensor_azimuth:long_name = "Sensor azimuth angle at pixel locations" ;
//		sensor_azimuth:units = "degrees" ;
//		sensor_azimuth:valid_min = -18000s ;
//		sensor_azimuth:valid_max = 18000s ;
//		sensor_azimuth:scale_factor = 0.01 ;
//		sensor_azimuth:add_offset = 0. ;
//	short sensor_zenith(number_of_scans, CCD_pixels) ;
//		sensor_zenith:_FillValue = -32767s ;
//		sensor_zenith:long_name = "Sensor zenith angle at pixel locations" ;
//		sensor_zenith:units = "degrees" ;
//		sensor_zenith:valid_min = 0s ;
//		sensor_zenith:valid_max = 18000s ;
//		sensor_zenith:scale_factor = 0.01 ;
//		sensor_zenith:add_offset = 0. ;
//	short solar_azimuth(number_of_scans, CCD_pixels) ;
//		solar_azimuth:_FillValue = -32767s ;
//		solar_azimuth:long_name = "Solar azimuth angle at pixel locations" ;
//		solar_azimuth:units = "degrees" ;
//		solar_azimuth:valid_min = -18000s ;
//		solar_azimuth:valid_max = 18000s ;
//		solar_azimuth:scale_factor = 0.01 ;
//		solar_azimuth:add_offset = 0. ;
//	short solar_zenith(number_of_scans, CCD_pixels) ;
//		solar_zenith:_FillValue = -32767s ;
//		solar_zenith:long_name = "Solar zenith angle at pixel locations" ;
//		solar_zenith:units = "degrees" ;
//		solar_zenith:valid_min = 0s ;
//		solar_zenith:valid_max = 18000s ;
//		solar_zenith:scale_factor = 0.01 ;
//		solar_zenith:add_offset = 0. ;
//	ubyte quality_flag(number_of_scans, CCD_pixels) ;
//		quality_flag:long_name = "Geolocation pixel quality flags" ;
//		quality_flag:flag_masks = 1UB, 2UB, 4UB ;
//		quality_flag:flag_meanings = "off_earth solar_eclipse terrain_bad" ;
//  } // group geolocation_data

group: navigation_data {
  variables:
  	float att_quat(number_of_scans, quaternion_elements) ;
  		att_quat:_FillValue = -32767.f ;
  		att_quat:long_name = "Attitude quaternions at EV mid-times" ;
  		att_quat:valid_min = -1.f ;
  		att_quat:valid_max = 1.f ;
  	float att_ang(number_of_scans, vector_elements) ;
  		att_ang:_FillValue = -32767.f ;
  		att_ang:long_name = "Attitude angles (roll, pitch, yaw) at EV mid-times" ;
  		att_ang:units = "degrees" ;
  		att_ang:valid_min = -180.f ;
  		att_ang:valid_max = 180.f ;
  	float orb_pos(number_of_scans, vector_elements) ;
  		orb_pos:_FillValue = -9999999.f ;
  		orb_pos:long_name = "Orbit position vectors at EV mid-times (ECR)" ;
  		orb_pos:units = "meters" ;
  		orb_pos:valid_min = -7100000.f ;
  		orb_pos:valid_max = 7100000.f ;
  	float orb_vel(number_of_scans, vector_elements) ;
  		orb_vel:_FillValue = -32767.f ;
  		orb_vel:long_name = "Orbit velocity vectors at EV mid-times (ECR)" ;
  		orb_vel:units = "meters/second" ;
  		orb_vel:valid_min = -7600.f ;
  		orb_vel:valid_max = 7600.f ;
  	float tilt_angle(number_of_scans) ;
  		tilt_angle:long_name = "OCI tilt angle at EV mid-times" ;
  		tilt_angle:units = "degrees" ;
  		tilt_angle:_FillValue = -32767.f ;
  		tilt_angle:valid_min = -22.5f ;
  		tilt_angle:valid_max = 20.5f ;
//  	float CCD_scan_angles(number_of_scans, CCD_pixels) ;
//  		CCD_scan_angles:long_name = "Scan angles for blue and red band science pixels" ;
//  		CCD_scan_angles:units = "degrees" ;
//  		CCD_scan_angles:_FillValue = -32767.f ;
//  		CCD_scan_angles:valid_min = -110.f ;
//  		CCD_scan_angles:valid_max = 250.f ;
//  	float SWIR_scan_angles(number_of_scans, SWIR_pixels) ;
//  		SWIR_scan_angles:long_name = "Scan angles for SWIR band science pixels" ;
//  		SWIR_scan_angles:units = "degrees" ;
//  		SWIR_scan_angles:_FillValue = -32767.f ;
//  		SWIR_scan_angles:valid_min = -110.f ;
//  		SWIR_scan_angles:valid_max = 250.f ;
  } // group navigation_data

group: observation_data {
  variables:
//  	float rhot_blue(blue_bands, number_of_scans, ccd_pixels) ;
//  		rhot_blue:_FillValue = -32767.f ;
//  		rhot_blue:long_name = "Top of Atmosphere Blue Band Reflectance" ;
//  		rhot_blue:valid_min = 0.f ;
//  		rhot_blue:valid_max = 1.3 ;
//  		rhot_blue:units = "dimensionless" ;
//  	byte qual_blue(blue_bands, number_of_scans, ccd_pixels) ;
//  		qual_blue:_FillValue = 255b ;
//  		qual_blue:long_name = "Blue Band Quality Flag" ;
//  		qual_blue:flag_masks = 1, 2, 4 ;
//  		qual_blue:flag_meanings = "saturation" ;
//  	float rhot_red(red_bands, number_of_scans, ccd_pixels) ;
//  		rhot_red:_FillValue = -32767.f ;
//  		rhot_red:long_name = "Top of Atmosphere Red Band Reflectance" ;
//  		rhot_red:valid_min = 0.f ;
//  		rhot_red:valid_max = 1.3 ;
//  		rhot_red:units = "dimensionless" ;
//  	byte qual_red(red_bands, number_of_scans, ccd_pixels) ;
//  		qual_red:_FillValue = 255b ;
//  		qual_red:long_name = "Red Band Quality Flag" ;
//  		qual_red:flag_masks = 1, 2, 4 ;
//  		qual_red:flag_meanings = "saturation" ;
//  	float rhot_SWIR(SWIR_bands, number_of_scans, ccd_pixels) ;
//  		rhot_SWIR:_FillValue = -32767.f ;
//  		rhot_SWIR:long_name = "Top of Atmosphere SWIR Band Reflectance" ;
//  		rhot_SWIR:valid_min = 0.f ;
//  		rhot_SWIR:valid_max = 1.3 ;
//  		rhot_SWIR:units = "dimensionless" ;
//  	byte qual_SWIR(SWIR_bands, number_of_scans, ccd_pixels) ;
//  		qual_SWIR:_FillValue = 255b ;
//  		qual_SWIR:long_name = "SWIR Band Quality Flag" ;
//  		qual_SWIR:flag_masks = 1, 2, 4 ;
//  		qual_SWIR:flag_meanings = "saturation" ;
  } // group observation_data
}
